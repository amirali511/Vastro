module vastro

// Solar constants
pub const solar_mass 							= 1.989e30 // kg
pub const solar_radius 						= 6.957e8 // m
pub const solar_apparent_magnitude = -26.74 // mag
pub const solar_luminosity	 				= 3.828e26 // W
pub const solar_absolute_magnitude = 4.83 // mag
pub const solar_temperature 				= 5778 // K

// Gravitational constants
pub const gravitational_constant 		= 6.67430e-11 // m^3 kg^-1 s^-2

// Light and wave constants
pub const speed_of_light 						= 3e8 // m/s
pub const boltzmann_constant 				= 1.380649e-23 // J/K
pub const stefan_boltzmann_constant 	= 5.670374419e-8 // W m^-2 K^-4
pub const plank_constant 						= 6.62607015e-34 // J s	
pub const planck_constant_reduced 		= 1.054571817e-34 // J s

// Distance constants
pub const au 												= 1.495978707e11 // m
pub const light_year 								= 9.4607304725808e15 // m
pub const parsec 										= 3.0856775814913673e16 // m

// Earth constants
pub const earth_mass = 5.972e24 // kg
pub const earth_radius = 6.371e6 // m
pub const earth_temperature = 288 // K
pub const earth_albedo = 0.306