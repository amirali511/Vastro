module vastro

// Solar constants
pub const solar_mass 							= 1.989e30 // kg
pub const solar_radius 						= 6.957e8 // m
pub const solar_apparent_magnitude = -26.74 // mag
pub const solar_luminosity	 				= 3.828e26 // W
pub const solar_absolute_magnitude = 4.83 // mag
pub const solar_temperature 				= 5778 // K